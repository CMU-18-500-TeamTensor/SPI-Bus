`default_nettype none

module ChipInterface ();



endmodule : ChipInterface